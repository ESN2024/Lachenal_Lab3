
module lab3_qs (
	clk_clk,
	reset_reset_n,
	opencores_i2c_0_export_0_scl_pad_io,
	opencores_i2c_0_export_0_sda_pad_io);	

	input		clk_clk;
	input		reset_reset_n;
	inout		opencores_i2c_0_export_0_scl_pad_io;
	inout		opencores_i2c_0_export_0_sda_pad_io;
endmodule
